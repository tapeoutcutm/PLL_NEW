VERSION 5.8 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO tt_um_Improved_delay_PLL
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 161000 BY 225760 ;
  SYMMETRY X Y ;

  ###########################################################
  # Power Pins
  ###########################################################
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0 224560 161000 225760 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0 0 161000 1200 ;
    END
  END VGND

  ###########################################################
  # Control Pins
  ###########################################################
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000 0 3000 2000 ;
    END
  END clk

  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4000 0 5000 2000 ;
    END
  END ena

  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6000 0 7000 2000 ;
    END
  END rst_n

  ###########################################################
  # ui_in[0..7]
  ###########################################################
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8000 0 9000 2000 ;
    END
  END ui_in[0]

  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10000 0 11000 2000 ;
    END
  END ui_in[1]

  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12000 0 13000 2000 ;
    END
  END ui_in[2]

  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14000 0 15000 2000 ;
    END
  END ui_in[3]

  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16000 0 17000 2000 ;
    END
  END ui_in[4]

  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18000 0 19000 2000 ;
    END
  END ui_in[5]

  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20000 0 21000 2000 ;
    END
  END ui_in[6]

  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22000 0 23000 2000 ;
    END
  END ui_in[7]

  ###########################################################
  # uo_out[0..7]
  ###########################################################
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000 223760 3000 225760 ;
    END
  END uo_out[0]

  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4000 223760 5000 225760 ;
    END
  END uo_out[1]

  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6000 223760 7000 225760 ;
    END
  END uo_out[2]

  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8000 223760 9000 225760 ;
    END
  END uo_out[3]

  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10000 223760 11000 225760 ;
    END
  END uo_out[4]

  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12000 223760 13000 225760 ;
    END
  END uo_out[5]

  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14000 223760 15000 225760 ;
    END
  END uo_out[6]

  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16000 223760 17000 225760 ;
    END
  END uo_out[7]

  ###########################################################
  # uio_in[0..7]
  ###########################################################
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24000 0 25000 2000 ;
    END
  END uio_in[0]

  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26000 0 27000 2000 ;
    END
  END uio_in[1]

  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28000 0 29000 2000 ;
    END
  END uio_in[2]

  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30000 0 31000 2000 ;
    END
  END uio_in[3]

  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32000 0 33000 2000 ;
    END
  END uio_in[4]

  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34000 0 35000 2000 ;
    END
  END uio_in[5]

  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36000 0 37000 2000 ;
    END
  END uio_in[6]

  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38000 0 39000 2000 ;
    END
  END uio_in[7]

  ###########################################################
  # uio_out[0..7]
  ###########################################################
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24000 223760 25000 225760 ;
    END
  END uio_out[0]

  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26000 223760 27000 225760 ;
    END
  END uio_out[1]

  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28000 223760 29000 225760 ;
    END
  END uio_out[2]

  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30000 223760 31000 225760 ;
    END
  END uio_out[3]

  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32000 223760 33000 225760 ;
    END
  END uio_out[4]

  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34000 223760 35000 225760 ;
    END
  END uio_out[5]

  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36000 223760 37000 225760 ;
    END
  END uio_out[6]

  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38000 223760 39000 225760 ;
    END
  END uio_out[7]

  ###########################################################
  # uio_oe[0..7]
  ###########################################################
  PIN uio_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24000 111880 25000 113880 ;
    END
  END uio_oe[0]

  PIN uio_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26000 111880 27000 113880 ;
    END
  END uio_oe[1]

  PIN uio_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28000 111880 29000 113880 ;
    END
  END uio_oe[2]

  PIN uio_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30000 111880 31000 113880 ;
    END
  END uio_oe[3]

  PIN uio_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32000 111880 33000 113880 ;
    END
  END uio_oe[4]

  PIN uio_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34000 111880 35000 113880 ;
    END
  END uio_oe[5]

  PIN uio_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36000 111880 37000 113880 ;
    END
  END uio_oe[6]

  PIN uio_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38000 111880 39000 113880 ;
    END
  END uio_oe[7]

END MACRO

END LIBRARY
