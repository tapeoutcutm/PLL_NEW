VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

SITE core
  CLASS CORE ;
  SIZE 1 BY 1 ;
  SYMMETRY X Y ;
END core

MACRO tt_um_Improved_delay_PLL
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 161.000 BY 225.760 ;
  SYMMETRY X Y ;
  SITE core ;

  # ---------------------------
  # Signal Pins
  # ---------------------------
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3000 0 4000 2000 ;
    END
  END clk

  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5000 0 6000 2000 ;
    END
  END ena

  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7000 0 8000 2000 ;
    END
  END rst_n

  # ui_in[0..7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9000 0 10000 2000 ;
    END
  END ui_in[0]

  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11000 0 12000 2000 ;
    END
  END ui_in[1]

  # ... repeat for ui_in[2..7]

  # uo_out[0..7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13000 225760 14000 227760 ;
    END
  END uo_out[0]

  # ... repeat for uo_out[1..7]

  # uio_in/out/oe[0..7] (bi-directional interface pins)
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15000 0 16000 2000 ;
    END
  END uio_in[0]

  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15000 225760 16000 227760 ;
    END
  END uio_out[0]

  PIN uio_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15000 10000 16000 12000 ;
    END
  END uio_oe[0]

  # ---------------------------
  # Power Pins
  # ---------------------------
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0 224560 161000 225760 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0 0 161000 1200 ;
    END
  END VGND

END tt_um_Improved_delay_PLL
END LIBRARY
