VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO PFD
  CLASS CORE ;
  FOREIGN PFD ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.670 BY 6.400 ;
  SITE unithddb1 ;
  PIN Clk_Ref
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.879000 ;
    ANTENNADIFFAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 2.420 5.520 3.520 5.710 ;
        RECT 2.420 5.210 2.650 5.520 ;
        RECT 0.040 1.740 0.310 3.510 ;
        RECT 0.040 1.450 2.100 1.740 ;
    END
  END Clk_Ref
  PIN Up
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.427200 ;
    PORT
      LAYER li1 ;
        RECT 6.270 4.780 6.560 5.780 ;
        RECT 6.390 4.040 6.560 4.780 ;
        RECT 6.260 3.560 6.560 4.040 ;
    END
  END Up
  PIN Down
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.427200 ;
    PORT
      LAYER li1 ;
        RECT 6.520 1.930 6.810 2.930 ;
        RECT 6.640 1.190 6.810 1.930 ;
        RECT 6.510 0.710 6.810 1.190 ;
    END
  END Down
  PIN Clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.879000 ;
    ANTENNADIFFAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 0.900 2.060 1.230 2.230 ;
        RECT 4.700 1.850 4.890 2.720 ;
        RECT 4.390 1.620 4.890 1.850 ;
      LAYER mcon ;
        RECT 0.980 2.060 1.150 2.230 ;
      LAYER met1 ;
        RECT 0.710 2.010 1.210 2.290 ;
    END
  END Clk2
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 4.340 3.290 5.010 4.100 ;
        RECT 5.780 3.360 6.000 3.880 ;
        RECT 5.560 3.290 6.230 3.360 ;
        RECT 4.340 3.120 7.670 3.290 ;
        RECT 0.780 2.760 0.990 2.780 ;
        RECT 0.700 2.590 1.060 2.760 ;
        RECT 0.780 2.510 0.990 2.590 ;
        RECT 1.730 0.920 1.910 1.280 ;
        RECT 6.030 0.700 6.250 1.030 ;
      LAYER mcon ;
        RECT 4.940 3.120 5.110 3.290 ;
        RECT 5.280 3.120 5.450 3.290 ;
        RECT 5.620 3.120 5.790 3.290 ;
        RECT 5.960 3.120 6.130 3.290 ;
        RECT 6.300 3.120 6.470 3.290 ;
        RECT 6.640 3.120 6.810 3.290 ;
        RECT 0.800 2.590 0.970 2.760 ;
        RECT 1.740 1.010 1.910 1.180 ;
        RECT 6.070 0.780 6.240 0.950 ;
      LAYER met1 ;
        RECT 0.000 2.960 7.670 3.440 ;
        RECT 0.740 2.530 1.040 2.960 ;
        RECT 2.280 1.240 2.520 2.960 ;
        RECT 1.680 0.950 2.520 1.240 ;
        RECT 5.600 1.010 5.870 2.960 ;
        RECT 5.600 0.720 6.270 1.010 ;
    END
  END GND
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.890 5.350 7.670 6.400 ;
        RECT 1.370 4.790 7.670 5.350 ;
        RECT 5.050 4.600 7.670 4.790 ;
      LAYER li1 ;
        RECT 0.000 6.050 7.670 6.220 ;
        RECT 1.650 5.720 2.070 6.050 ;
        RECT 1.510 5.510 2.220 5.720 ;
        RECT 5.770 5.080 6.000 6.050 ;
      LAYER mcon ;
        RECT 0.800 6.050 0.970 6.220 ;
        RECT 1.140 6.050 1.310 6.220 ;
        RECT 1.480 6.050 1.650 6.220 ;
        RECT 1.820 6.050 1.990 6.220 ;
        RECT 2.160 6.050 2.330 6.220 ;
        RECT 2.500 6.050 2.670 6.220 ;
        RECT 2.840 6.050 3.010 6.220 ;
        RECT 3.180 6.050 3.350 6.220 ;
        RECT 3.520 6.050 3.690 6.220 ;
        RECT 3.860 6.050 4.030 6.220 ;
        RECT 4.200 6.050 4.370 6.220 ;
        RECT 4.540 6.050 4.710 6.220 ;
        RECT 4.880 6.050 5.050 6.220 ;
        RECT 5.220 6.050 5.390 6.220 ;
        RECT 5.560 6.050 5.730 6.220 ;
        RECT 5.900 6.050 6.070 6.220 ;
        RECT 6.240 6.050 6.410 6.220 ;
        RECT 6.580 6.050 6.750 6.220 ;
      LAYER met1 ;
        RECT 0.000 5.920 7.670 6.400 ;
    END
    PORT
      LAYER nwell ;
        RECT 6.770 3.070 7.670 3.080 ;
        RECT 4.430 2.950 7.670 3.070 ;
        RECT 3.970 1.570 7.670 2.950 ;
        RECT 3.970 0.310 5.140 1.570 ;
      LAYER li1 ;
        RECT 6.020 2.540 6.250 2.930 ;
        RECT 7.040 2.660 7.450 2.830 ;
        RECT 6.020 2.250 6.330 2.540 ;
        RECT 7.100 2.370 7.400 2.660 ;
        RECT 6.020 2.230 6.250 2.250 ;
        RECT 7.040 2.200 7.450 2.370 ;
        RECT 7.100 1.930 7.400 2.200 ;
        RECT 7.040 1.760 7.450 1.930 ;
        RECT 4.690 0.310 4.900 1.420 ;
        RECT 0.000 0.140 7.670 0.310 ;
      LAYER mcon ;
        RECT 6.160 2.310 6.330 2.480 ;
        RECT 7.140 2.180 7.350 2.390 ;
        RECT 0.800 0.140 0.970 0.310 ;
        RECT 1.140 0.140 1.310 0.310 ;
        RECT 1.480 0.140 1.650 0.310 ;
        RECT 1.820 0.140 1.990 0.310 ;
        RECT 2.160 0.140 2.330 0.310 ;
        RECT 2.500 0.140 2.670 0.310 ;
        RECT 2.840 0.140 3.010 0.310 ;
        RECT 3.180 0.140 3.350 0.310 ;
        RECT 3.520 0.140 3.690 0.310 ;
        RECT 3.860 0.140 4.030 0.310 ;
        RECT 4.200 0.140 4.370 0.310 ;
        RECT 4.540 0.140 4.710 0.310 ;
        RECT 4.880 0.140 5.050 0.310 ;
        RECT 5.220 0.140 5.390 0.310 ;
        RECT 5.560 0.140 5.730 0.310 ;
        RECT 5.900 0.140 6.070 0.310 ;
        RECT 6.240 0.140 6.410 0.310 ;
        RECT 6.580 0.140 6.750 0.310 ;
      LAYER met1 ;
        RECT 6.100 2.250 7.410 2.540 ;
        RECT 6.560 2.070 7.410 2.250 ;
        RECT 6.560 0.480 6.860 2.070 ;
        RECT 0.000 0.000 7.670 0.480 ;
    END
  END VDPWR
  OBS
      LAYER li1 ;
        RECT 1.550 4.880 2.240 5.240 ;
        RECT 0.370 4.630 2.240 4.880 ;
        RECT 2.840 5.040 3.550 5.230 ;
        RECT 0.370 3.950 0.640 4.630 ;
        RECT 2.840 4.570 3.280 5.040 ;
        RECT 5.260 4.910 5.480 5.780 ;
        RECT 5.260 4.740 6.100 4.910 ;
        RECT 5.900 4.610 6.100 4.740 ;
        RECT 2.840 4.450 5.710 4.570 ;
        RECT 0.870 4.400 5.710 4.450 ;
        RECT 0.870 4.190 3.290 4.400 ;
        RECT 5.900 4.270 6.130 4.610 ;
        RECT 5.900 4.230 6.090 4.270 ;
        RECT 5.250 4.060 6.090 4.230 ;
        RECT 0.370 3.710 3.100 3.950 ;
        RECT 5.250 3.680 5.470 4.060 ;
        RECT 2.860 0.860 3.050 3.320 ;
        RECT 3.340 2.510 3.530 3.320 ;
        RECT 4.220 2.620 4.410 2.750 ;
        RECT 3.950 2.510 4.410 2.620 ;
        RECT 3.340 2.260 4.410 2.510 ;
        RECT 3.340 2.200 3.640 2.260 ;
        RECT 3.340 1.090 3.600 2.200 ;
        RECT 3.950 2.180 4.410 2.260 ;
        RECT 4.220 2.070 4.410 2.180 ;
        RECT 5.510 2.060 5.730 2.930 ;
        RECT 5.510 1.890 6.350 2.060 ;
        RECT 6.160 1.760 6.350 1.890 ;
        RECT 5.140 1.550 5.960 1.720 ;
        RECT 6.160 1.470 6.380 1.760 ;
        RECT 3.340 0.860 3.530 1.090 ;
        RECT 3.960 0.750 4.420 1.440 ;
        RECT 6.150 1.420 6.380 1.470 ;
        RECT 6.150 1.380 6.330 1.420 ;
        RECT 5.500 1.210 6.330 1.380 ;
        RECT 5.500 0.830 5.720 1.210 ;
      LAYER mcon ;
        RECT 2.870 1.240 3.040 1.410 ;
        RECT 3.430 2.230 3.600 2.400 ;
        RECT 5.200 1.550 5.370 1.720 ;
        RECT 4.090 1.000 4.260 1.170 ;
      LAYER met1 ;
        RECT 3.340 2.140 3.690 2.490 ;
        RECT 5.130 1.470 5.450 1.790 ;
        RECT 2.810 1.230 3.790 1.470 ;
        RECT 2.810 1.180 4.320 1.230 ;
        RECT 3.560 0.940 4.320 1.180 ;
      LAYER via ;
        RECT 3.370 2.170 3.660 2.460 ;
        RECT 5.160 1.500 5.420 1.760 ;
      LAYER met2 ;
        RECT 3.340 2.460 3.690 2.490 ;
        RECT 3.340 2.190 5.400 2.460 ;
        RECT 3.340 2.140 3.690 2.190 ;
        RECT 5.140 1.790 5.400 2.190 ;
        RECT 5.130 1.470 5.450 1.790 ;
  END
END PFD
END LIBRARY

